library verilog;
use verilog.vl_types.all;
entity bin_bcd_original_vlg_vec_tst is
end bin_bcd_original_vlg_vec_tst;
