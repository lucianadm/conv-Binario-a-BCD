library verilog;
use verilog.vl_types.all;
entity bin_3bcd_vlg_vec_tst is
end bin_3bcd_vlg_vec_tst;
